* NGSPICE file created from counter.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VNB VPB VGND VPWR A X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VPB VNB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VPB VNB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR A X VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 Q CLK D VPB VNB VPWR VGND
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_2 Q CLK D VPB VNB VPWR VGND
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X11 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X18 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X19 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X20 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X21 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X22 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X25 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_4 VGND VPWR VNB VPB Q D CLK
X0 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X1 a_1020_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X2 a_572_47# a_193_47# a_475_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X3 VPWR a_1062_300# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0913 ps=0.855 w=0.42 l=0.15
X4 a_634_183# a_475_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.149 ps=1.22 w=0.64 l=0.15
X5 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.109 ps=1.36 w=0.42 l=0.15
X7 a_475_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X8 VGND a_1062_300# a_1020_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X9 VPWR a_634_183# a_568_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X11 a_568_413# a_27_47# a_475_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0662 ps=0.735 w=0.42 l=0.15
X12 a_634_183# a_475_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X13 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0913 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_183# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X16 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.106 ps=0.975 w=0.65 l=0.15
X17 VGND a_891_413# a_1062_300# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X18 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X24 VPWR a_891_413# a_1062_300# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.28 ps=2.56 w=1 l=0.15
X25 a_891_413# a_193_47# a_634_183# VNB sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X26 a_475_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X27 VGND a_634_183# a_572_47# VNB sky130_fd_pr__nfet_01v8 ad=0.149 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X29 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 VPB VNB VGND VPWR A1 A2 B1 X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B X C VGND VPWR VPB VNB
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_1 VPWR VGND VPB VNB B1_N Y A1 A2
X0 a_300_297# a_27_413# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X3 Y a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.102 ps=0.99 w=0.65 l=0.15
X4 VPWR A1 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_384_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X6 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.111 ps=1.37 w=0.42 l=0.15
X7 a_300_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VPB VNB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 VGND VPWR A X VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 VNB VPB VPWR VGND A X B
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt counter VGND VPWR clk_i cnt_o[0] cnt_o[1] cnt_o[2] rst_n_i
XFILLER_0_94_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_76_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_73_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_95_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_69_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_66_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_4_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_73_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_387 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_75_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Right_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_64_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Right_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_77_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_79_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_75_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Right_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_89_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_99_Left_201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_77_Right_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_91_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Right_86 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_99_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_95_Right_95 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_73_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_18_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_74_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Left_147 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_61_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_71_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_54_Left_156 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_79_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_19_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_87_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Left_174 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_Left_183 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_90_Left_192 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_93_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_101_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_16_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_85_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_89_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_99_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_67_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_86_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_75_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_100_Left_202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_68_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_74_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_101_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_75_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_86_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_79_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_10_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_101_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_69_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_57_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_79_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_95_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_48_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Left_180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_85_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_98_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_77_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Right_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_67_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_67_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Right_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_59_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_80_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_82_Right_82 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_91_Right_91 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_83_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_86_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_65_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_116 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_68_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_83_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Left_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_87_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_87_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Left_143 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Left_152 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_97_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_69_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_79_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f_clk_i VGND VPWR VGND VPWR clknet_0_clk_i clknet_1_0__leaf_clk_i sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_108 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_82_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Left_199 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_86_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_18_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_97_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_87_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09_ VGND VPWR _00_ _07_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_1_Right_1 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_98_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_98_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_73_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_73_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_97_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_97_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_66_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_69_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_522 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_40_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_79_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_79_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08_ _07_ net2 net1 VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_95_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_87_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_140 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_66_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_69_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_68_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_95_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Right_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_98_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_42_Right_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_98_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Right_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_77_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_95_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_95_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_99_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_76_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Right_89 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_98_Right_98 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_81_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_94_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_66_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_66_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_2_Left_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_98_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_98_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Left_168 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_77_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_85_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Left_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_72_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_84_Left_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_95_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Left_195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_64_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_73_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_46_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_85_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_67_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_96_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_96_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_70_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_76_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_78_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_21_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_89_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_96_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_98_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_71_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_98_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_66_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_66_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_85_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_46_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_96_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_70_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_78_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_58_Right_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_78_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Right_67 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_98_Left_200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Right_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Right_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Right_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_57_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_76_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_89_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Left_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_97_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Left_146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Left_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_76_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_62_Left_164 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_32_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Left_173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Left_182 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk_i VGND VPWR VGND VPWR clk_i clknet_0_clk_i sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_46_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_83_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 VGND VPWR rst_n_i net1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_93_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_97_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_8_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_75_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_8_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_79_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_79_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_82_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_19_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_6_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_83_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_96_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_78_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_75_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_75_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_94_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_97_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_79_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_86_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_69_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Left_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_170 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_32_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Right_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_93_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_46_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_46_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_100_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_96_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Right_63 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_75_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Right_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_Right_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_90_Right_90 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_62_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_384 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_94_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_94_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_13_Left_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_95_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Left_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_76_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_99_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_40_Left_142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_94_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_58_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_95_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_107 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_100_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_87_Left_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_96_Left_198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_62_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_38_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_75_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_396 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_94_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_73_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_44_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_94_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_73_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_89_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_73_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_87_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_98_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_66_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_89_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_36_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_76_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_92_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_60_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_87_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_95_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_87_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Right_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_87_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Right_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_95_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_50_Right_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_59_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_101_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_99_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_95_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_4_Right_4 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_81_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Right_79 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Right_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Right_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_58_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_37_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_87_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_87_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_95_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_79_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_56_Left_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_74_Left_176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_69_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_85_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_69_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_61_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_92_Left_194 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_58_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_88_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_89_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_92_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_67_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_79_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_43_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_100_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Left_191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_67_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_57_Right_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_66_Right_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_86_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Right_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_84_Right_84 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_82_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_93_Right_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_99_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_99_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_2_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_89_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_16_Left_118 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_86_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_55_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_136 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_97_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Left_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_92_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Left_154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Left_172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_74_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_79_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_98_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_75_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_86_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_86_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_73_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_412 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_101_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_96_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Right_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_59_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_83_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_34_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_69_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18_ net4 clknet_1_1__leaf_clk_i _02_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_16_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_98_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Left_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_55_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_72_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Right_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_98_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_35_Right_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_54_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_77_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Right_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Right_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_91_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Right_80 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_98_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_73_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_86_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_55_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Left_123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_68_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_30_Left_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_83_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_62_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_11_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_85_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17_ net3 clknet_1_0__leaf_clk_i _01_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_94_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_101_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_98_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_98_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_66_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_72_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Left_179 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_95_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Left_188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Left_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_98_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_78_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_83_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_78_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16_ VGND VPWR VGND VPWR net2 _00_ clknet_1_0__leaf_clk_i sky130_fd_sc_hd__dfxtp_4
XFILLER_0_87_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_61_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_66_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_85_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_77_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_46_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_96_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_7_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_73_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_84_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15_ VPWR VGND VGND VPWR _05_ _06_ net1 _02_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_66_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_89_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_48_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_71_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_66_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_85_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_85_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Right_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_53_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Right_40 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_98_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_99_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_77_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_49_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_58_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Right_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_52_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_12_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Right_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14_ net4 net3 _06_ net2 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_87_Right_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_34_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_96_Right_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_96_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_8_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Left_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Left_139 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_46_Left_148 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_55_Left_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_98_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_64_Left_166 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_82_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Left_175 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_93_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Left_184 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_77_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_Left_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_96_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_96_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_387 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_43_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13_ VPWR VGND VPWR VGND net4 _05_ net2 net3 sky130_fd_sc_hd__a21boi_1
XFILLER_0_75_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_45_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_97_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_101_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_56_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Left_203 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_58_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_95_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_95_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_67_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_77_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_85_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_96_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_67_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_96_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12_ VGND VPWR _01_ _04_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_38_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_78_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_101_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_79_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_94_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_409 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_94_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_56_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_68_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Left_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_64_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_88_Left_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_80_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_clk_i VGND VPWR VGND VPWR clknet_0_clk_i clknet_1_1__leaf_clk_i sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_96_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_96_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Right_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11_ VPWR VGND _04_ _03_ net1 VPWR VGND sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_47_Right_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_75_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_56_Right_56 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_65_Right_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_91_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_78_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Right_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_62_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Right_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_92_Right_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_57_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_96_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_100_Right_100 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_89_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_76_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_126 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_79_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_135 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Left_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_89_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput2 VGND VPWR net2 cnt_o[0] VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_82_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_80_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_64_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10_ VGND VPWR VPWR VGND net2 _03_ net3 sky130_fd_sc_hd__xor2_1
XFILLER_0_83_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_83_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_94_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_31_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_76_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_99_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_79_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_50_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_89_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_89_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_97_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 net1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_21_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_87_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_79_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xoutput3 VPWR VGND cnt_o[1] net3 VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_50_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_78_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_78_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_51_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_83_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_94_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_73_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_2 net2 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_21_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_76_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_76_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_94_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_94_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput4 VGND VPWR net4 cnt_o[2] VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Left_150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_58_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_66_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_16_Right_16 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_87_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_25_Right_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Right_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_59_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_43_Right_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_61_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_69_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Right_61 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_80_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_88_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_67_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_96_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Right_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_78_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_94_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_59_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Left_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_53_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_76_Left_178 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Left_187 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_56_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_101_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Left_196 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_7_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_88_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_4_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_67_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_81_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_94_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
.ends

