* NGSPICE file created from counter.ext - technology: sky130A

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VNB VPB VGND VPWR A X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VPB VNB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VPB VNB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR A X VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 X A VPB VNB VGND VPWR
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 Q CLK D VPB VNB VPWR VGND
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_2 Q CLK D VPB VNB VPWR VGND
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X11 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X18 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X19 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X20 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X21 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X22 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X25 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR X B A C VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_1 VPWR VGND VPB VNB A2 A1 B1 X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_1 VPB VNB VGND VPWR A B Y C
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND VPB VNB A2 A1 B1 Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 VGND VPWR A X VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 B1 Y A1 VPB VNB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt counter VGND VPWR clk_i cnt_o[0] cnt_o[1] cnt_o[2] rst_n_i
XFILLER_0_27_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_48_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_58_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_58_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_52_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_56_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_153 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_62_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_30_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_53_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_84 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Right_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_49_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Right_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_19_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Left_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Left_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_49_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_19_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_23_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_34_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_39_Left_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Left_112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_54_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_54_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_42_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_46_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_27_Left_91 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_57_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_11_Left_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_Right_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_54_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_9 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_46_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_clk_i VGND VPWR VGND VPWR clknet_0_clk_i clknet_1_0__leaf_clk_i sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09_ VGND VPWR _00_ _07_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_1_Right_1 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08_ _07_ net2 net1 VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_11_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_79 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_48_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Right_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Right_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_54_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_48_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_82 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Left_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Left_118 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_59_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_67 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_58_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_46_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_63_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_50_Left_114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_23_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_58_Right_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_48_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk_i VGND VPWR VGND VPWR clk_i clknet_0_clk_i sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_23_Left_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_62_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xinput1 VGND VPWR rst_n_i net1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_26_Left_90 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Left_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_61_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Left_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_63_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Right_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Right_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_61_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Right_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Right_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Right_54 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Right_63 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_315 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_62_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_327 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_44_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_58_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_58_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_32_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_95 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_58_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Right_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Right_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Left_108 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_53_Left_117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_126 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Right_4 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_35_Left_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Left_123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_49_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_10_Right_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_86 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Left_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1 net5 net3 VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Right_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Right_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 net6 _01_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Left_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Left_110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18_ net4 clknet_1_1__leaf_clk_i _02_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Left_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Right_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_53_Right_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Right_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_54_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_80 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_58_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_62_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17_ net3 clknet_1_0__leaf_clk_i net6 VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_58_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_30_Left_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_47_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16_ net2 clknet_1_0__leaf_clk_i _00_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_47_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15_ VGND VPWR _02_ _06_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_48_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Right_40 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_43_Left_107 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_52_Left_116 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_49_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14_ VGND VPWR _06_ _04_ net1 _05_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_34_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_98 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_21_Left_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13_ VPWR VGND VPWR VGND net3 net2 net4 _05_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_45_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_56_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12_ VPWR VGND VGND VPWR net2 net3 _04_ net4 sky130_fd_sc_hd__nand3_1
XFILLER_0_7_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_46_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Left_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_52_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_39_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_clk_i VGND VPWR VGND VPWR clknet_0_clk_i clknet_1_1__leaf_clk_i sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_29_Right_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_56_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11_ VPWR VGND VPWR VGND net5 net2 _03_ _01_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_47_Right_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Right_56 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_28_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xoutput2 VGND VPWR net2 cnt_o[0] VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10_ VGND VPWR net5 net1 _03_ net2 VPWR VGND sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_25_Left_89 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_28_Left_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_12_Left_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput3 VGND VPWR net3 cnt_o[1] VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_64 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_100 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_166 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput4 VGND VPWR net4 cnt_o[2] VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_58_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Right_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_34_Right_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_43_Right_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_52_Right_52 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_61_Right_61 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_55_Left_119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Right_2 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
.ends

